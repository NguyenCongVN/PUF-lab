`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 03/25/2017 01:55:31 PM
// Design Name:
// Module Name: dflipflop
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////


module dflipflop(input D,
                 input Clk,
                 output reg Q);
    always @ (posedge Clk) begin
        Q <= D;
    end
endmodule
