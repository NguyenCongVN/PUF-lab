or  O1(D, SA, SB);


module lut_or (
    output reg D,
    input wire SA,
    input wire SB
);
    
endmodule